package ascii;

    typedef enum logic [7:0] 
    {
        // numbers
        ZERO = 8'h30,
        ONE = 8'h31,
        TWO = 8'h32,
        THREE = 8'h33,
        FOUR = 8'h34,
        FIVE = 8'h35,
        SIX = 8'h36,
        SEVEN = 8'h37, 
        EIGHT = 8'h38,
        NINE = 8'h39,

        // Uppercase Letters
        CHAR_A_U = 8'h41,
        CHAR_B_U = 8'h42,
        CHAR_C_U = 8'h43,
        CHAR_D_U = 8'h44,
        CHAR_E_U = 8'h45,
        CHAR_F_U = 8'h46,
        CHAR_G_U = 8'h47,
        CHAR_H_U = 8'h48,
        CHAR_I_U = 8'h49,
        CHAR_J_U = 8'h4A,
        CHAR_K_U = 8'h4B,
        CHAR_L_U = 8'h4C,
        CHAR_M_U = 8'h4D,
        CHAR_N_U = 8'h4E,
        CHAR_O_U = 8'h4F,
        CHAR_P_U = 8'h50,
        CHAR_Q_U = 8'h51,
        CHAR_R_U = 8'h52,
        CHAR_S_U = 8'h53,
        CHAR_T_U = 8'h54,
        CHAR_U_U = 8'h55,
        CHAR_V_U = 8'h56,
        CHAR_W_U = 8'h57,
        CHAR_X_U = 8'h58,
        CHAR_Y_U = 8'h59,
        CHAR_Z_U = 8'h5A,
    
        // Lowercase Letters
        CHAR_A_L = 8'h61,
        CHAR_B_L = 8'h62,
        CHAR_C_L = 8'h63,
        CHAR_D_L = 8'h64,
        CHAR_E_L = 8'h65,
        CHAR_F_L = 8'h66,
        CHAR_G_L = 8'h67,
        CHAR_H_L = 8'h68,
        CHAR_I_L = 8'h69,
        CHAR_J_L = 8'h6A,
        CHAR_K_L = 8'h6B,
        CHAR_L_L = 8'h6C,
        CHAR_M_L = 8'h6D,
        CHAR_N_L = 8'h6E,
        CHAR_O_L = 8'h6F,
        CHAR_P_L = 8'h70,
        CHAR_Q_L = 8'h71,
        CHAR_R_L = 8'h72,
        CHAR_S_L = 8'h73,
        CHAR_T_L = 8'h74,
        CHAR_U_L = 8'h75,
        CHAR_V_L = 8'h76,
        CHAR_W_L = 8'h77,
        CHAR_X_L = 8'h78,
        CHAR_Y_L = 8'h79,
        CHAR_Z_L = 8'h7A,

        // Other Characters
        COLON = 8'h3A,
        STOP = 8'h2E,
        SEMI_COLON = 8'h3B,
        MINUS = 8'h2D,
        DIVIDE = 8'h2F,
        PLUS = 8'h2B,
        COMMA = 8'h2C,
        LESS_THAN = 8'h3C,
        GREATER_THAN = 8'h3E,
        EQUALS = 8'h3D,
        QUESTION = 8'h3F,
        DOLLAR = 8'h24,
        SPACE = 8'h20,
        EXCLAIM = 8'h21

    } e_character;

endpackage